
            .out_cnt(out_cnt),
            .rx_dac_gain(rx_dac_gain),
            .is_10_bit(is_10_bit),
            .adc_clk_dly(adc_clk_dly),
            .ld_dac_en(ld_dac_en),
            .ld_dac_val(ld_dac_val),
            .adc_chb_result(adc_chb_result),
            .adc_cha_result(adc_cha_result),
            .adc_fco_result(adc_fco_result),
            .adc_dco_result(adc_dco_result),
            .adc_spi_wr_en(adc_spi_wr_en),
            .adc_spi_rd_en(adc_spi_rd_en),
            .adc_spi_busy(adc_spi_busy),
            .adc_spi_wdata(adc_spi_wdata),
            .adc_spi_wr_len(adc_spi_wr_len),
            .adc_spi_rdata(adc_spi_rdata),
            .rx_dac_spi_wr_en(rx_dac_spi_wr_en),
            .rx_dac_spi_busy(rx_dac_spi_busy),
            .rx_dac_spi_wdata(rx_dac_spi_wdata),
            .l_adc_spi_rd_en(l_adc_spi_rd_en),
            .l_adc_spi_busy(l_adc_spi_busy),
            .l_adc_spi_rdata1(l_adc_spi_rdata1),
            .l_adc_spi_rdata(l_adc_spi_rdata),
            .timer_l(timer_l),
            .timer_rst(timer_rst),
            .timer_stop(timer_stop),
            .timer_h(timer_h),