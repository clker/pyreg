
            .spi_rw_len(spi_rw_len),
            .spi_rcv_rise_align(spi_rcv_rise_align),
            .spi_busy(spi_busy),
            .spi_ch_sel(spi_ch_sel),
            .spi_send_rise_align(spi_send_rise_align),
            .out_cnt(out_cnt),
            .rx_dac_gain(rx_dac_gain),
            .is_10_bit(is_10_bit),
            .adc_clk_dly(adc_clk_dly),
            .spi_wdata(spi_wdata),
            .spi_wr_en(spi_wr_en),
            .spi_rd_en(spi_rd_en),
            .adc_fifo_rd_en(adc_fifo_rd_en),
            .adc_fifo_rst(adc_fifo_rst),
            .ld_dac_en(ld_dac_en),
            .ld_dac_val(ld_dac_val),
            .adc_fifo_empty(adc_fifo_empty),
            .adc_fifo_full(adc_fifo_full),
            .adc_chb_result(adc_chb_result),
            .adc_cha_result(adc_cha_result),
            .adc_fco_result(adc_fco_result),
            .adc_dco_result(adc_dco_result),
            .spi_rdata1(spi_rdata1),
            .spi_rdata(spi_rdata),